RMS value calculation of a file.

*
V1 N1 0 AC 1V SIN(0V 1V 1KHz)
R1 N1 0 1k

.ac dec 10 1Hz 1KHz

.tran 0.01ms 1ms

.END
